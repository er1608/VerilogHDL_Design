library verilog;
use verilog.vl_types.all;
entity edge_dff_vlg_vec_tst is
end edge_dff_vlg_vec_tst;
