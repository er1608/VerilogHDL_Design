`timescale 1ns/100ps
module Testbench();
	reg[2:0] A, B;
	reg Cin;
	wire[3:0] S, mS;
	
	initial
	begin
		#640 $stop;
	end
	
	initial
	begin
		Gen();
	end
	
	Adder Inst1(.A(A), .B(B), .Cin(Cin), .S(S));
	//CLA_M Inst2 (.A(A), .B(B), .Cin(Cin), .S(mS));
	
	task Gen;
	begin
		A<=0;
		B<=0;
		Cin<=0;
		forever begin
		#5 A <= (A + 1);
			if (A == 3'b111)
			begin
				#0 B <= (B + 1);
				if (B == 3'b111)
				begin
					#0 Cin <= (Cin+1);
				end
			end
			if ((S==mS))
				#0 $display ("Expected result: %d .Simulation result: %d --> PASS",S ,mS);
			else	
				#0	$display ("Expected result: %d .Simulation result: %d --> FAIL",S ,mS);
			end
		end
	endtask
endmodule
