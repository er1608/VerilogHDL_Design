library verilog;
use verilog.vl_types.all;
entity AU2_pipeline_vlg_vec_tst is
end AU2_pipeline_vlg_vec_tst;
